DC Power Supply with a BJT Series Regulator
*Rohan Rajesh Kalbag - 20D170033

.model bc547a NPN IS=10f BF=200 ISE=10.3f IKF=50m NE=1.3 
+ BR=9.5 VAF=80 IKR=12m ISC=47p NC=2 VAR=10 RB=280 RE=1 RC=40 
+ tr=0.3u tf=0.5n cje=12p vje=0.48 mje=0.5 cjc=6p vjc=0.7 mjc=0.33 kf=2f 
 
.model SL100 NPN IS=100f BF=80 ISE=10.3f IKF=50m NE=1.3 
+ BR=9.5 VAF=80 IKR=12m ISC=47p NC=2 VAR=10 RB=100 RE=1 RC=10 
+ tr=0.3u tf=0.5n cje=12p vje=0.48 mje=0.5 cjc=6p vjc=0.7 mjc=0.33 kf=2f

.SUBCKT ZENER_12 1 2
D1 1 2 DF
DZ 3 1 DR
VZ 2 3 4.4
.MODEL DF D(IS =27.5p RS=0.620 N=1.10 CJO =78.3p VJ=1.00 M =0.330 TT =50.1n)
.MODEL DR D(IS =5.49f RS=50 N=1.77 )
.ENDS

v1 1 0 dc
rc 1 2 1k
q1 1 2 3 SL100
q2 2 4 5 bc547a
x1 0 5 ZENER_12
r1 3 4 10.21k
r2 4 0 14.79k
rl 3 0 1k

.dc v1 15 25 0.5
.control
run
plot v(3) vs v(1)
.endc
.end