Question 1
*Rohan Rajesh Kalbag - 20D170033

.include TL084.txt

v1 3 0 dc 15
v2 4 0 dc -15
x1 1 2 3 4 5 TL084
vi 6 0 0.1 ac
r1 6 1 6.8k
l1 1 0 1

.ac dec 10 10m 10k
.control
run
plot vdb(5) - vdb(6) xlog
.endc
.end