Photo Diode - Rohan Rajesh Kalbag - 20d170033

.include lm324.txt
v1 3 0 ac 0 dc 5 
r2 2 5 13.7k
r3 2 0 280
x1 2 1 3 0 5 lm324
c2 2 0 1u
r1 1 5 1.4Meg
c1 1 5 3.3p
vref 2 0 dc 0.1 ac 0
i1 1 0 ac 0 dc 
cj 1 0 11p

.dc i1 0 2.4u 0.1u
.control
run
plot v(5)
.endc
.end
