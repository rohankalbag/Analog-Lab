RC Integrator
*Components
r1 1 2 10k
c1 2 0 0.1u
*pulse of width 0.00001s = 0.01RC, height 1, and period 0.00002s
V1 1 0 pulse(0 1 0 0 0 0.00001 0.00002)
*Analysis Command
.tran 0.000001 0.00006
.control 
run
plot v(1) v(2)
.endc
.end