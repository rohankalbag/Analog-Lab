Full Wave Precision Rectifier
*Rohan Rajesh Kalbag - 20D170033

.include ua741.txt
.include Diode_1N914.txt

v1 2 0 dc 15
v2 3 0 dc -15
vi 5 0 sin(0 5 1k 0 0 0)

*half-wave-precision-rectifier

.subckt HWPR 1 2 3 4 5 6 7
x1 1 2 3 4 5 ua741
d1 5 2 1N914
d2 7 5 1N914
r1 6 2 10k
r2 2 7 10k
.include ua741.txt
.include Diode_1N914.txt
.ends

*inverting summer
x3 0 1 2 3 4 5 6 HWPR
r3 5 8 10k
r4 6 8 5k
x2 0 8 2 3 9 ua741
r5 8 9 10k
rl 9 0 1k

.tran 1ms 10ms
.control
run
plot v(9) v(5)
.endc
.end