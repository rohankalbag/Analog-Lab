Midsem Q2d
*Rohan Rajesh Kalbag - 20D170033

.include lm324.txt

v1 3 0 dc 5
v2 4 0 dc -5
x1 1 8 3 4 5 lm324
vin 2 0 dc
vos 7 8 dc 0.002
vref 6 0 dc 1.2235 ac 0
r1 6 1 9.5k 
r2 1 0 10.1k
rg 2 7 3.234k
rf 7 5 57.68k 
.control
dc vin 0 2 1m
plot v(5)
.endc
.end