Inverting Amplifier with Opamp-2
*Rohan Rajesh Kalbag - 20D170033

.include ua741.txt

v1 2 0 dc 15
v2 3 0 dc -15
x1 0 1 2 3 4 ua741
vi 5 0 sin(0 2 1k 0 0 0)
r1 5 1 1k
r2 1 4 10k

.tran 1ms 10ms
.control
run
plot v(5) v(4)
.endc
.end