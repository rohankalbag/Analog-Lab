RC lowpass filter
*Components
r1 1 2 10k
c1 2 0 0.1u
V1 1 0 dc 0 ac 1 $ac analysis
*Analysis Command
.ac dec 10 1 10k 
.control 
run
plot vdb(2)
.endc
.end