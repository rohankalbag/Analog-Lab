Unregulated DC supply without capacitive filter

.include Diode_1N914.txt
r 3 4 1k
d1 1 3 1N914
d2 4 1 1N914
d3 2 3 1N914
d4 4 2 1N914
v1 1 2 sin(0 21.213 50 0 0 0)

.tran v1 0.02m 60m

.control

run
plot v(3)-v(4)

.endc
.end
