RC Differentiator
*Components
c1 1 2 0.1u
r1 2 0 10k
V1 1 0 pulse(0 5 0 0 0 10m 20m)
*Analysis Command
.tran 0.02m 60m
.control 
run
plot v(1) v(2)
.endc
.end