RC circuit transient analysis

*describe circuit
*<element-name> <nodes> <value/model>
r1 1 2 1k
r2 2 0 1k
v 1 0 pwl(0 0 10m 0 11m 5 20m 5)

*analysis command
.tran 10u 20ms
.control

run

*display command
plot v(1) v(2)
.endc 

.end
