RC Integrator
*Components
r1 1 2 10k
c1 2 0 0.1u
V1 1 0 pulse(0 5 0 0 0 0.0001 0.0002)
*Analysis Command
.tran 0.0001m 0.0006
.control 
run
plot v(1) v(2)
.endc
.end