RC bandpass filter

*Components
r1 1 2 10k
c1 2 3 0.1u
r2 3 0 10k
c2 3 0 0.1u
V1 1 0 dc 0 ac 1 $ac analysis

*Analysis Command
.ac dec 500 1m 10Meg 
.control 
run
plot vdb(3)
print vdb(3)
.endc
.end

