Single Pole Active High Pass Filter 
*Rohan Rajesh Kalbag 20D170033
.include "ua741.txt"
*after calculating theoretical f_c = (1/(2pi*R*C)) = 338.62Hz
*we see -3dB frequency as ~ f_c 

x1 1 2 3 4 5 ua741
v1 3 0 12 dc
v2 4 0 -12 dc
r1 5 2 9.1k
r2 2 0 1k
ra 1 0 4.7k
ca 6 1 0.1u
vi 6 0 dc 0 ac 1
.ac dec 10 10m 100Meg
.control
run
plot vdb(5)-vdb(6) xlog
plot {57.29*(vp(5)-vp(6))} xlog
.endc
.end