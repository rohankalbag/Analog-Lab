RLC bandpass filter

*Components
l1 1 2 10m
c1 2 3 0.1u
r2 3 0 1k
V1 1 0 dc 0 ac 1 $ac analysis

*Analysis Command
.ac dec 10 10m 1000Meg 
.control 
run
plot vdb(3)
.endc
.end

