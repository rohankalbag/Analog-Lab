RC Differentiator
*Components
c1 1 2 0.1u
r1 2 0 10k
V1 1 0 pulse(0 5 0 0 0 0.001 0.002)
*Analysis Command
.tran 0.002m 0.006
.control 
run
plot v(1) v(2)
.endc
.end