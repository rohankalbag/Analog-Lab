RC circuit transient analysis

*describe circuit
*<element-name> <nodes> <value/model>
r1 1 2 1k
c 2 0 1u
v 1 0 sin(0 2 1k 0 0)

*analysis command
.tran 10u 20ms
.control

run

*display command
plot v(1) v(2)
.endc 

.end
