Inverting Amplifier with Opamp
*Rohan Rajesh Kalbag - 20D170033

.include ua741.txt

v1 2 0 dc 15
v2 3 0 dc -15
x1 0 1 2 3 4 ua741
vi 5 0 0.1 ac
r1 5 1 1k
r2 1 4 10k

.ac dec 10 10m 10Meg
.control
run
plot vdb(4) - vdb(5)
print vdb(4) - vdb(5)
.endc
.end