Full Wave Precision Rectifier
*Rohan Rajesh Kalbag - 20D170033

.include ua741.txt
.include Diode_1N914.txt

*half-wave-rectifier
v1 2 0 dc 15
v2 3 0 dc -15
x1 0 1 2 3 4 ua741
d1 4 1 1N914
d2 6 4 1N914
vi 5 0 sin(0 5 1k 0 0 0)
r1 5 1 10k
r2 1 6 10k

*inverting summer
r3 5 8 10k
r4 6 8 5k
x2 0 8 2 3 9 ua741
r5 8 9 10k
rl 9 0 1k

.tran 1ms 10ms
.control
run
plot v(9) v(5)
.endc
.end