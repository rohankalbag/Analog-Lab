OPAMP based circuit - 3 
*Rohan Rajesh Kalbag - 20D170033

.include ua741.txt

.SUBCKT ZENER_12 1 2
D1 1 2 DF
DZ 3 1 DR
VZ 2 3 3.5
.MODEL DF D(IS =27.5p RS=0.620 N=1.10 CJO =78.3p VJ=1.00 M =0.330 TT =50.1n)
.MODEL DR D(IS =5.49f RS=50 N=1.77 )
.ENDS

v1 2 0 dc 15
v2 3 0 dc -15
x1 1 0 2 3 4 ua741
r1 8 1 8.2k
r2 1 6 15k
r3 4 6 1k
x2 6 7 ZENER_12
x3 0 7 ZENER_12
x4 0 9 2 3 8 ua741
r4 6 9 18k
c1 9 8 47n
r5 9 8 1.5Meg

.tran 10us 101ms 99ms
.control
run
plot v(8) v(6)
.endc
.end