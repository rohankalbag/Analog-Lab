RC Integrator
*Components
r1 1 2 10k
c1 2 0 0.1u
V1 1 0 pulse(0 5 0 0 0 0.001 0.002)
*Analysis Command
.tran 0.001m 0.006
.control 
run
plot v(1) v(2)
.endc
.end