OPAMP based circuit - 3 
*Rohan Rajesh Kalbag - 20D170033

.include ua741.txt

v1 2 0 dc 15
v2 3 0 dc -15
x1 0 1 2 3 4 ua741
vi 5 0 pulse(2 -2 0 0 0 0.5ms 1ms 0)
r1 5 1 18k
c1 1 4 47n
r2 1 4 1.5Meg
.tran 10us 110ms 100ms
.control
run
plot v(4)
.endc
.end