Photo Diode Bode Plot
*Rohan Rajesh Kalbag - 20d170033

.include lm324.txt
v1 3 0 dc 5 
r2 2 5 13.7k
r3 2 0 280
x1 2 1 3 0 5 lm324
c2 2 0 1u
r1 1 5 1.4Meg
c1 1 5 3.3p
vref 2 0 0.1
i1 1 6 dc 1.5u ac
vd 6 0 0 
cj 1 0 11p

.ac dec 10 10 100Meg
.control
run
plot {20*log(abs(v(5)/i(vd)))} xlog
.endc
.end
