OPAMP based circuit - 1
*Rohan Rajesh Kalbag - 20D170033

.include lm324.txt

v1 3 0 dc 5
c1 3 0 0.01u
x1 1 2 3 0 5 lm324
vi 1 0 dc
rl 5 0 10k
rf 2 5 180k
rg 6 5 20k
c2 6 0 0.01u
r1 3 6 75k
r2 6 0 820

.dc vi 0.1 5 0.1
.control
run
plot v(5) v(1)
plot v(5) vs v(1)
.endc
.end